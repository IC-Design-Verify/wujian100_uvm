`ifdef USE_ADDR_MAP
  `include "addr_map/tb_addr_map_pre_module.v"
`endif
`ifdef USE_HAD
  `include "had/tb_had_pre_module.v"
`endif
//module top_sim();
//
//endmodule
