`ifndef TOP_SIM_TESTCASE_PACKAGE__SV
`define TOP_SIM_TESTCASE_PACKAGE__SV
`include "soc_subsys_top_sim_seq_pkg.svh"

//package top_sim_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "subsys_top_sim_testcase.svh"

  //import addr_map_testcase_pkg::*;
  //import had_testcase_pkg::*;

//endpackage

`include "addr_map/addr_map_testcase_pkg.svh"
`include "had/had_testcase_pkg.svh"

`endif
