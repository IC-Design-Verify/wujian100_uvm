`ifdef USE_APB0_WDT
  `include "apb0_wdt/tb_apb0_wdt_post_module.v"
`endif
`ifdef USE_APB0_PWM
  `include "apb0_pwm/tb_apb0_pwm_post_module.v"
`endif
`ifdef USE_APB0_USI
  `include "apb0_usi/tb_apb0_usi_post_module.v"
`endif
//module apb0();
//
//endmodule
