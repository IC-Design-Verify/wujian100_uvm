//interface assignment

// Sub Environment Interface assignment 

