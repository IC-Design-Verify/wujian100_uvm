`ifndef AHB_HS_TESTCASE_PACKAGE__SV
`define AHB_HS_TESTCASE_PACKAGE__SV
`include "soc_subsys_ahb_hs_seq_pkg.svh"

//package ahb_hs_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "subsys_ahb_hs_testcase.svh"

  //import soc_dma_testcase_pkg::*;

//endpackage

`include "soc_dma/soc_dma_testcase_pkg.svh"

`endif
