`ifndef GATE_SIM_TESTCASE_PACKAGE__SV
`define GATE_SIM_TESTCASE_PACKAGE__SV
`include "soc_subsys_gate_sim_seq_pkg.svh"

//package gate_sim_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "subsys_gate_sim_testcase.svh"

  //import sdf_sim_testcase_pkg::*;

//endpackage

`include "sdf_sim/sdf_sim_testcase_pkg.svh"

`endif
