`ifndef AHB_LS_TESTCASE_PACKAGE__SV
`define AHB_LS_TESTCASE_PACKAGE__SV
`include "soc_subsys_ahb_ls_seq_pkg.svh"

//package ahb_ls_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;
  import ahb_pkg::*;


  
  //
  `include "subsys_ahb_ls_testcase.svh"


//endpackage


`endif
