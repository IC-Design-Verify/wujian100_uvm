//module apb0_usi();
//
//endmodule
