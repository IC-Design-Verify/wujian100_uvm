`ifndef SOC_SUBSYS_HAD_SEQ_PKG__SV
`define SOC_SUBSYS_HAD_SEQ_PKG__SV
//package soc_subsys_had_seq_pkg;
  //import uvm_pkg::*;
  //import soc_top_vseq_lib_pkg::*;
  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;

  `include "soc_top_v_sequence_pkg.svh"
  `include "soc_subsys_top_sim_seq_pkg.svh"

  //
  `include "had/soc_had_sequence.svh"
  `include "had/soc_had_vseq.svh"

//endpackage
`endif
