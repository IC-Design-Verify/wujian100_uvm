//module sdf_sim();
//
//endmodule
