`ifndef SOC_TOP_V_SEQUENCE_PACKAGE__SV
`define SOC_TOP_V_SEQUENCE_PACKAGE__SV

  //vip package

  //vip package, sub_env needs

  //agent package

  //reg_model package

  //env package
  import soc_top_env_pkg::*;

  //sub_env sequence_pkg

  //include reg_sequence

  //include intr_sequence

  `include "soc_top_v_sequence_base.svh"
  //include v_sequence
  `include "soc_top_v_sequence.svh"

  //include other sequences

`endif
