`ifndef SDF_SIM_TESTCASE_PACKAGE__SV
`define SDF_SIM_TESTCASE_PACKAGE__SV
`include "sdf_sim/soc_sdf_sim_seq_pkg.svh"

//package sdf_sim_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "sdf_sim/sdf_sim_testcase.svh"


//endpackage


`endif
