//module soc_dma();
//
//endmodule
