//module ahb_ls();
//
//endmodule
