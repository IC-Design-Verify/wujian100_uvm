//module apb1_pmu();
//
//endmodule
