`ifdef USE_SOC_DMA
  `include "soc_dma/tb_soc_dma_pre_module.v"
`endif
//module ahb_hs();
//
//endmodule
