`ifndef SOC_TOP_TESTCASE__SV
`define SOC_TOP_TESTCASE__SV

  //vip package

  

  //reg_model package

  //m_env package
  //import soc_top_env_pkg::*;

  //import soc_top_intr_seq_pkg::*;
  //reg_seq package

  //include test_base
  `include "soc_top_test_base.svh"

  //include testcase
  `include "soc_top_test_lib.svh"

`endif
