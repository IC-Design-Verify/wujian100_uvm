`ifndef APB0_PWM_TESTCASE_PACKAGE__SV
`define APB0_PWM_TESTCASE_PACKAGE__SV
`include "apb0_pwm/soc_apb0_pwm_seq_pkg.svh"

//package apb0_pwm_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "apb0_pwm/apb0_pwm_testcase.svh"


//endpackage


`endif
