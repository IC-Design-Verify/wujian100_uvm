//module had();
//
//endmodule
