`ifndef SOC_TOP_INTR_SEQ_PACKAGE__SV
`define SOC_TOP_INTR_SEQ_PACKAGE__SV
package soc_top_intr_sequence_pkg;
  import uvm_pkg::*;

  //agent package

  //reg_model package

  //env package
  import soc_top_env_pkg::*;

  // include intr_sequence
  `include "soc_top_intr_sequence_base.svh"

endpackage
`endif
