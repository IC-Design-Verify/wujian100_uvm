`ifndef APB1_RTC_TESTCASE_PACKAGE__SV
`define APB1_RTC_TESTCASE_PACKAGE__SV
`include "apb1_rtc/soc_apb1_rtc_seq_pkg.svh"

//package apb1_rtc_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "apb1_rtc/apb1_rtc_testcase.svh"


//endpackage


`endif
