`ifndef HAD_TESTCASE_PACKAGE__SV
`define HAD_TESTCASE_PACKAGE__SV
`include "had/soc_had_seq_pkg.svh"

//package had_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "had/had_testcase.svh"


//endpackage


`endif
