`ifndef SOC_DMA_TESTCASE_PACKAGE__SV
`define SOC_DMA_TESTCASE_PACKAGE__SV
`include "soc_dma/soc_soc_dma_seq_pkg.svh"

//package soc_dma_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "soc_dma/soc_dma_testcase.svh"


//endpackage


`endif
