`ifndef ADDR_MAP_TESTCASE_PACKAGE__SV
`define ADDR_MAP_TESTCASE_PACKAGE__SV
`include "addr_map/soc_addr_map_seq_pkg.svh"

//package addr_map_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;
  import ahb_pkg::*;


  
  //
  `include "addr_map/addr_map_testcase.svh"


//endpackage


`endif
