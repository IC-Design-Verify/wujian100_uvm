//module addr_map();
//
//endmodule
