`ifndef APB1_GPIO_TESTCASE_PACKAGE__SV
`define APB1_GPIO_TESTCASE_PACKAGE__SV
`include "apb1_gpio/soc_apb1_gpio_seq_pkg.svh"

//package apb1_gpio_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;
  import ahb_pkg::*;


  
  //
  `include "apb1_gpio/apb1_gpio_testcase.svh"


//endpackage


`endif
