`ifndef APB0_USI_TESTCASE_PACKAGE__SV
`define APB0_USI_TESTCASE_PACKAGE__SV
`include "apb0_usi/soc_apb0_usi_seq_pkg.svh"

//package apb0_usi_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;


  
  //
  `include "apb0_usi/apb0_usi_testcase.svh"


//endpackage


`endif
