//module apb0_wdt();
//
//endmodule
