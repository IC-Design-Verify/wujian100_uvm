`ifndef SOC_TOP_DEFINE__SV
`define SOC_TOP_DEFINE__SV

    `define MERGE_ITF_NAME(prename, name) prename``name
    `define HIER_SOC_TOP tb_top.dut

    //-----------------------------------------------------------
    //-----------------------------------------------------------

    //Sub Env Define

`endif
