//module apb1_gpio();
//
//endmodule
