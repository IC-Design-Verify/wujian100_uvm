//module apb1_rtc();
//
//endmodule
