//module apb0_pwm();
//
//endmodule
