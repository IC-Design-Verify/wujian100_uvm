`ifndef APB1_PMU_TESTCASE_PACKAGE__SV
`define APB1_PMU_TESTCASE_PACKAGE__SV
`include "apb1_pmu/soc_apb1_pmu_seq_pkg.svh"

//package apb1_pmu_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;
  import ahb_pkg::*;


  
  //
  `include "apb1_pmu/apb1_pmu_testcase.svh"


//endpackage


`endif
