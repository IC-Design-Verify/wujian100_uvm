`ifdef USE_APB1_RTC
  `include "apb1_rtc/tb_apb1_rtc_post_module.v"
`endif
`ifdef USE_APB1_GPIO
  `include "apb1_gpio/tb_apb1_gpio_post_module.v"
`endif
`ifdef USE_APB1_PMU
  `include "apb1_pmu/tb_apb1_pmu_post_module.v"
`endif
//module apb1();
//
//endmodule
