`ifndef APB0_WDT_TESTCASE_PACKAGE__SV
`define APB0_WDT_TESTCASE_PACKAGE__SV
`include "apb0_wdt/soc_apb0_wdt_seq_pkg.svh"

//package apb0_wdt_testcase_pkg;
  //import uvm_pkg::*;

  //import svt_uvm_pkg::*;
  //import svt_ahb_uvm_pkg::*;    
  //import svt_ahb_sequence_pkg::*;
  import ahb_pkg::*;


  
  //
  `include "apb0_wdt/apb0_wdt_testcase.svh"


//endpackage


`endif
