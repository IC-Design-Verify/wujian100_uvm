`ifdef USE_SDF_SIM
  `include "sdf_sim/tb_sdf_sim_post_module.v"
`endif
//module gate_sim();
//
//endmodule
