`ifndef SOC_TOP_TESTS__SV
`define SOC_TOP_TESTS__SV

`include "soc_top_v_sequence_pkg.svh"
`include "soc_top_testcase_pkg.svh"
  `include "subsys_apb0_testcase_pkg.svh"
  `include "subsys_apb1_testcase_pkg.svh"
  `include "subsys_gate_sim_testcase_pkg.svh"
  `include "subsys_ahb_hs_testcase_pkg.svh"
  `include "subsys_ahb_ls_testcase_pkg.svh"
  `include "subsys_top_sim_testcase_pkg.svh"


`endif
